library verilog;
use verilog.vl_types.all;
entity break_sv is
end break_sv;
